`define ADDR_WIDTH 10
`define DATA_WIDTH 32
